/*
Authors: Krzysztof Korbaś, Emilia Jerdanek
*/

import snake_pkg::*;

module mode_control(
    input logic clk,

    output wire game_mode mode
);

endmodule 
