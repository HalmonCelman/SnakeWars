/*
Authors: Krzysztof Korbaś, Emilia Jerdanek
*/

package snake_pkg;

typedef enum { 
    MENU,
    ERROR,
    GAME,
    ENDSCR
} game_mode;

endpackage