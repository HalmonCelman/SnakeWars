/*
Authors: Krzysztof Korbaś, Emilia Jerdanek
*/
`timescale 1 ns / 1 ps

import snake_pkg::*;

module top (
    input  wire clk100MHz,
    input  wire clk,
    input  wire rst,
    input  wire rx,
    
    output logic tx,
    output logic hsync,
    output logic vsync,
    output logic [RGB_B-1:0] rgb,

    inout wire mouse_clk,
    inout wire mouse_data
);

map_s map, map_nxt;
vga_if vga_in(), vga_out();
logic [11:0] mouse_x, mouse_y;
direction dir_int, dir2_int;
logic clk_divided;
logic left_int, right_int;
logic rcvdir;
logic eaten1, eaten2;

assign hsync = vga_out.hsync;
assign vsync = vga_out.vsync;

vga_timing u_vga_timing(
    .clk,
    .rst,
    .vga(vga_in)
);

draw u_draw (
    .clk,
    .rst,
    .map,
    .mouse_x,
    .mouse_y,
    .mode(GAME),
    .vga_in,
    .vga_out,
    .rgb
);

clk_div u_clk_div(
    .clk,
    .rst,
    .clk_divided
);

collisons u_collisions(
    .map,
    .map_nxt,
    .mode(GAME),
    
    .eaten1,
    .eaten2,
    .won(),
    .lost(),
    .draw()
);

move u_move (
    .clk,
    .clk_div(clk_divided),
    .rst,
    .dir1(dir_int),
    .dir2(dir2_int),
    .rcvdir,
    .map,
    .predicted_map(map_nxt),
    .com_err(),
    .eaten1,
    .eaten2
);

mouse_move u_mouse_move (
    .clk,
    .clk_divided,
    .rst,
    .left(left_int),
    .right(right_int),
    .dir(dir_int)
);

mouse_control u_mouse_control(
    .clk100MHz,
    .clk75MHz(clk),
    .rst,
    .left(left_int),
    .right(right_int),
    .ps2_clk(mouse_clk),
    .ps2_data(mouse_data),
    .x(mouse_x),
    .y(mouse_y)
);

communicate u_communicate(
    .clk,
    .rst,
    .rx,
    .send(clk_divided),
    .tx,
    .dir1(dir_int),
    .dir2(dir2_int),
    .rcvdir
);

endmodule
